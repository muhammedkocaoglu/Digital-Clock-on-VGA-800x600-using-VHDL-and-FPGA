library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity vga800x600 is
	port(
		CLOCK_50		: in std_logic;
		KEY         : in std_logic_vector(2 downto 0);
		SW 			: in std_logic_vector(1 downto 0);
		rst         : in std_logic;  --key[3]
		
		--Outputs
		GPIO_0      : out std_logic_vector(1 downto 0);  --gpio[0] is for buzzer. 
		TD_RESET 	: out std_logic:='1';
		LEDR        : out std_logic_vector(1 downto 0);
		VGA_CLK     : out std_logic;
		VGA_BLANK   : out std_logic;
		VGA_HS,VGA_VS : inout std_logic;
		VGA_R,VGA_G,VGA_B : out std_logic_vector(9 downto 0)
	);
end entity;


architecture vga800x600 of vga800x600 is
	signal reset: std_logic:='0';
	signal clk_40: std_logic;
	signal clk_1hz: std_logic;
	signal cntr59: integer:=0; 
	signal cntr59_min: integer:=0;
	signal cntr59_hour: integer:=0;
	signal clk_div : std_logic_vector(20 downto 0);
	signal clk15 : std_logic;
	signal enable : std_logic;

----------------------------------------------------------------
   component PLL is
        port (
            clk_in_clk  : in  std_logic := 'X'; -- clk
            reset_reset : in  std_logic := 'X'; -- reset
            clk_out_clk : out std_logic         -- clk
        );
    end component PLL;
----------------------------------------------------------------
	constant HD : integer := 799;         --  639   Horizontal Display (640)
	constant HFP : integer := 40;         --   16   Right border (front porch)
	constant HSP : integer := 128;        --   96   Sync pulse (Retrace)
	constant HBP : integer := 88;         --   48   Left boarder (back porch)
	
	constant VD : integer := 599;         --  479   Vertical Display (480)
	constant VFP : integer := 1;       	  --   10   Right border (front porch)
	constant VSP : integer := 4;			  --    2   Sync pulse (Retrace)
	constant VBP : integer := 23;         --   33   Left boarder (back porch)
	
	signal hPos : integer := 0;
	signal vPos : integer := 0;
	
	signal videoOn : std_logic := '0';
	
		--Hafıza
	type HFZ is array (0 to 79) of std_logic_vector(0 to 39);
								
		constant BM_0: HFZ :=("0000000000000000000000000000000000000000",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0111000000000000000000000000000000001110",--5
									 "0111000000000000000000000000000000001110",--6
									 "0111000000000000000000000000000000001110",--7
									 "0111000000000000000000000000000000001110",--8
									 "0111000000000000000000000000000000001110",--9
								    "0111000000000000000000000000000000001110",--10         --0
								    "0111000000000000000000000000000000001110",--11
								    "0111000000000000000000000000000000001110",--12
								    "0111000000000000000000000000000000001110",--13
								    "0111000000000000000000000000000000001110",--14
								    "0111000000000000000000000000000000001110",--15
								    "0111000000000000000000000000000000001110",--16
								    "0111000000000000000000000000000000001110",--17
								    "0111000000000000000000000000000000001110",--18
								    "0111000000000000000000000000000000001110",--19
								    "0111000000000000000000000000000000001110",     --20
									 "0111000000000000000000000000000000001110",--1
								    "0111000000000000000000000000000000001110",--2
								    "0111000000000000000000000000000000001110",--3
								    "0111000000000000000000000000000000001110",--4
									 "0111000000000000000000000000000000001110",--5
									 "0111000000000000000000000000000000001110",--6
									 "0111000000000000000000000000000000001110",--7
									 "0111000000000000000000000000000000001110",--8
									 "0111000000000000000000000000000000001110",--9
								    "0111000000000000000000000000000000001110",--10         --0
								    "0111000000000000000000000000000000001110",--11
								    "0111000000000000000000000000000000001110",--12
								    "0111000000000000000000000000000000001110",--13
								    "0111000000000000000000000000000000001110",--14
								    "0111000000000000000000000000000000001110",--15
								    "0111000000000000000000000000000000001110",--16
								    "0111000000000000000000000000000000001110",--17
								    "0111000000000000000000000000000000001110",--18
								    "0111000000000000000000000000000000001110",--19
								    "0111000000000000000000000000000000001110",     --40
									 "0111000000000000000000000000000000001110",--1
								    "0111000000000000000000000000000000001110",--2
								    "0111000000000000000000000000000000001110",--3
								    "0111000000000000000000000000000000001110",--4
									 "0111000000000000000000000000000000001110",--5
									 "0111000000000000000000000000000000001110",--6
									 "0111000000000000000000000000000000001110",--7
									 "0111000000000000000000000000000000001110",--8
									 "0111000000000000000000000000000000001110",--9
								    "0111000000000000000000000000000000001110",--10         --0
								    "0111000000000000000000000000000000001110",--11
								    "0111000000000000000000000000000000001110",--12
								    "0111000000000000000000000000000000001110",--13
								    "0111000000000000000000000000000000001110",--14
								    "0111000000000000000000000000000000001110",--15
								    "0111000000000000000000000000000000001110",--16
								    "0111000000000000000000000000000000001110",--17
								    "0111000000000000000000000000000000001110",--18
								    "0111000000000000000000000000000000001110",--19
								    "0111000000000000000000000000000000001110",    --60
									 "0111000000000000000000000000000000001110",--1
								    "0111000000000000000000000000000000001110",--2
								    "0111000000000000000000000000000000001110",--3
								    "0111000000000000000000000000000000001110",--4
									 "0111000000000000000000000000000000001110",--5
									 "0111000000000000000000000000000000001110",--6
									 "0111000000000000000000000000000000001110",--7
									 "0111000000000000000000000000000000001110",--8
									 "0111000000000000000000000000000000001110",--9
								    "0111000000000000000000000000000000001110",--10         --0
								    "0111000000000000000000000000000000001110",--11
								    "0111000000000000000000000000000000001110",--12
								    "0111000000000000000000000000000000001110",--13
								    "0111000000000000000000000000000000001110",--14
								    "0111000000000000000000000000000000001110",--15
								    "0111000000000000000000000000000000001110",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0000000000000000000000000000000000000000");  --80
									 
	   constant BM_BOS:HFZ:=("0000000000000000000000000000000000000000",--1
								    "0000000000000000000000000000000000000000",--2
								    "0000000000000000000000000000000000000000",--3
								    "0000000000000000000000000000000000000000",--4
									 "0000000000000000000000000000000000000000",--5
									 "0000000000000000000000000000000000000000",--6
									 "0000000000000000000000000000000000000000",--7
									 "0000000000000000000000000000000000000000",--8
									 "0000000000000000000000000000000000000000",--9
								    "0000000000000000000000000000000000000000",--10         --BOS
								    "0000000000000000000000000000000000000000",--11
								    "0000000000000000000000000000000000000000",--12
								    "0000000000000000000000000000000000000000",--13
								    "0000000000000000000000000000000000000000",--14
								    "0000000000000000000000000000000000000000",--15
								    "0000000000000000000000000000000000000000",--16
								    "0000000000000000000000000000000000000000",--17
								    "0000000000000000000000000000000000000000",--18
								    "0000000000000000000000000000000000000000",--19
								    "0000000000000000000000000000000000000000",     --20
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000");
									 
										 
									 
									 
	   constant BM_1:HFZ:=  ("0000000000000000000000000000000000000000",--1
								    "0000000000000000000000000000000000001110",--2
								    "0000000000000000000000000000000000001110",--3
								    "0000000000000000000000000000000000001110",--4
									 "0000000000000000000000000000000000001110",--5
									 "0000000000000000000000000000000000001110",--6
									 "0000000000000000000000000000000000001110",--7
									 "0000000000000000000000000000000000001110",--8
									 "0000000000000000000000000000000000001110",--9
								    "0000000000000000000000000000000000001110",--10         --1
								    "0000000000000000000000000000000000001110",--11
								    "0000000000000000000000000000000000001110",--12
								    "0000000000000000000000000000000000001110",--13
								    "0000000000000000000000000000000000001110",--14
								    "0000000000000000000000000000000000001110",--15
								    "0000000000000000000000000000000000001110",--16
								    "0000000000000000000000000000000000001110",--17
								    "0000000000000000000000000000000000001110",--18
								    "0000000000000000000000000000000000001110",--19
								    "0000000000000000000000000000000000001110",     --20
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000001110",
									 "0000000000000000000000000000000000000000");	
									 
	  constant BM_2: HFZ :=("0000000000000000000000000000000000000000",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0111111111111111111111111111111111111110",--5
									 "0000000000000000000000000000000000011110",--6
									 "0000000000000000000000000000000000011110",--7
									 "0000000000000000000000000000000000011110",--8
									 "0000000000000000000000000000000000011110",--9
								    "0000000000000000000000000000000000011110",--10         --22222222222
								    "0000000000000000000000000000000000011110",--11                  --222222222222
								    "0000000000000000000000000000000000011110",--12
								    "0000000000000000000000000000000000011110",--13
								    "0000000000000000000000000000000000011110",--14
								    "0000000000000000000000000000000000011110",--15
								    "0000000000000000000000000000000000011110",--16
								    "0000000000000000000000000000000000011110",--17
								    "0000000000000000000000000000000000011110",--18
								    "0000000000000000000000000000000000011110",--19
								    "0000000000000000000000000000000000011110",     --20
									 "0000000000000000000000000000000000011110",--1
								    "0000000000000000000000000000000000011110",--2
								    "0000000000000000000000000000000000011110",--3
								    "0000000000000000000000000000000000011110",--4
									 "0000000000000000000000000000000000011110",--5
									 "0000000000000000000000000000000000011110",--6
									 "0000000000000000000000000000000000011110",--7
									 "0000000000000000000000000000000000011110",--8
									 "0000000000000000000000000000000000011110",--9
								    "0000000000000000000000000000000000011110",--10         
								    "0000000000000000000000000000000000011110",--11
								    "0000000000000000000000000000000000011110",--12
								    "0000000000000000000000000000000000011110",--13
								    "0000000000000000000000000000000000011110",--14
								    "0000000000000000000000000000000000011110",--15
								    "0000000000000000000000000000000000011110",--16
								    "0000000000000000000000000000000000011110",--17
								    "0000000000000000000000000000000000011110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0111111111111111111111111111111111111110",     --40
									 "0111111111111111111111111111111111111110",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111100000000000000000000000000000000000",--3
								    "0111100000000000000000000000000000000000",--4
									 "0111100000000000000000000000000000000000",--5
									 "0111100000000000000000000000000000000000",--6
									 "0111100000000000000000000000000000000000",--7
									 "0111100000000000000000000000000000000000",--8
									 "0111100000000000000000000000000000000000",--9
								    "0111100000000000000000000000000000000000",--10         
								    "0111100000000000000000000000000000000000",--11
								    "0111100000000000000000000000000000000000",--12
								    "0111100000000000000000000000000000000000",--13
								    "0111100000000000000000000000000000000000",--14
								    "0111100000000000000000000000000000000000",--15
								    "0111100000000000000000000000000000000000",--16
								    "0111100000000000000000000000000000000000",--17
								    "0111100000000000000000000000000000000000",--18
								    "0111100000000000000000000000000000000000",--19
								    "0111100000000000000000000000000000000000",    --60
									 "0111100000000000000000000000000000000000",--1
								    "0111100000000000000000000000000000000000",--2
								    "0111100000000000000000000000000000000000",--3
								    "0111100000000000000000000000000000000000",--4
									 "0111100000000000000000000000000000000000",--5
									 "0111100000000000000000000000000000000000",--6
									 "0111100000000000000000000000000000000000",--7
									 "0111100000000000000000000000000000000000",--8
									 "0111100000000000000000000000000000000000",--9
								    "0111100000000000000000000000000000000000",--10         
								    "0111100000000000000000000000000000000000",--11
								    "0111100000000000000000000000000000000000",--12
								    "0111100000000000000000000000000000000000",--13
								    "0111100000000000000000000000000000000000",--14
								    "0111100000000000000000000000000000000000",--15
								    "0111111111111111111111111111111111111110",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0000000000000000000000000000000000000000");  --80

		  constant BM_3: HFZ :=("0000000000000000000000000000000000000000",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0111111111111111111111111111111111111110",--5
									 "0000000000000000000000000000000000011110",--6
									 "0000000000000000000000000000000000011110",--7
									 "0000000000000000000000000000000000011110",--8
									 "0000000000000000000000000000000000011110",--9
								    "0000000000000000000000000000000000011110",--10         --33333333
								    "0000000000000000000000000000000000011110",--11                
								    "0000000000000000000000000000000000011110",--12
								    "0000000000000000000000000000000000011110",--13
								    "0000000000000000000000000000000000011110",--14
								    "0000000000000000000000000000000000011110",--15
								    "0000000000000000000000000000000000011110",--16
								    "0000000000000000000000000000000000011110",--17
								    "0000000000000000000000000000000000011110",--18
								    "0000000000000000000000000000000000011110",--19
								    "0000000000000000000000000000000000011110",     --20
									 "0000000000000000000000000000000000011110",--1
								    "0000000000000000000000000000000000011110",--2
								    "0000000000000000000000000000000000011110",--3
								    "0000000000000000000000000000000000011110",--4
									 "0000000000000000000000000000000000011110",--5
									 "0000000000000000000000000000000000011110",--6
									 "0000000000000000000000000000000000011110",--7
									 "0000000000000000000000000000000000011110",--8
									 "0000000000000000000000000000000000011110",--9
								    "0000000000000000000000000000000000011110",--10         
								    "0000000000000000000000000000000000011110",--11
								    "0000000000000000000000000000000000011110",--12
								    "0000000000000000000000000000000000011110",--13
								    "0000000000000000000000000000000000011110",--14
								    "0000000000000000000000000000000000011110",--15
								    "0000000000000000000000000000000000011110",--16
								    "0000000000000000000000000000000000011110",--17
								    "0000000000000000000000000000000000011110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0111111111111111111111111111111111111110",     --40
									 "0111111111111111111111111111111111111110",--1
								    "0111111111111111111111111111111111111110",--2
								    "0000000000000000000000000000000000011110",--3
								    "0000000000000000000000000000000000011110",--4
									 "0000000000000000000000000000000000011110",--5
									 "0000000000000000000000000000000000011110",--6
									 "0000000000000000000000000000000000011110",--7
									 "0000000000000000000000000000000000011110",--8
									 "0000000000000000000000000000000000011110",--9
								    "0000000000000000000000000000000000011110",--10         
								    "0000000000000000000000000000000000011110",--11
								    "0000000000000000000000000000000000011110",--12
								    "0000000000000000000000000000000000011110",--13
								    "0000000000000000000000000000000000011110",--14
								    "0000000000000000000000000000000000011110",--15
								    "0000000000000000000000000000000000011110",--16
								    "0000000000000000000000000000000000011110",--17
								    "0000000000000000000000000000000000011110",--18
								    "0000000000000000000000000000000000011110",--19
								    "0000000000000000000000000000000000011110",    --60
									 "0000000000000000000000000000000000011110",--1
								    "0000000000000000000000000000000000011110",--2
								    "0000000000000000000000000000000000011110",--3
								    "0000000000000000000000000000000000011110",--4
									 "0000000000000000000000000000000000011110",--5
									 "0000000000000000000000000000000000011110",--6
									 "0000000000000000000000000000000000011110",--7
									 "0000000000000000000000000000000000011110",--8
									 "0000000000000000000000000000000000011110",--9
								    "0000000000000000000000000000000000011110",--10         
								    "0000000000000000000000000000000000011110",--11
								    "0000000000000000000000000000000000011110",--12
								    "0000000000000000000000000000000000011110",--13
								    "0000000000000000000000000000000000011110",--14
								    "0000000000000000000000000000000000011110",--15
								    "0111111111111111111111111111111111111110",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0000000000000000000000000000000000000000");  --80
									 
		
		constant BM_4: HFZ :=("0000000000000000000000000000000000000000",--1
								    "0111100000000000000000000000000000011110",--2
								    "0111100000000000000000000000000000011110",--3
								    "0111100000000000000000000000000000011110",--4
									 "0111100000000000000000000000000000011110",--5
									 "0111100000000000000000000000000000011110",--6
									 "0111100000000000000000000000000000011110",--7
									 "0111100000000000000000000000000000011110",--8
									 "0111100000000000000000000000000000011110",--9
								    "0111100000000000000000000000000000011110",--10         --33333333
								    "0111100000000000000000000000000000011110",--11                
								    "0111100000000000000000000000000000011110",--12
								    "0111100000000000000000000000000000011110",--13
								    "0111100000000000000000000000000000011110",--14
								    "0111100000000000000000000000000000011110",--15
								    "0111100000000000000000000000000000011110",--16
								    "0111100000000000000000000000000000011110",--17
								    "0111100000000000000000000000000000011110",--18
								    "0111100000000000000000000000000000011110",--19
								    "0111100000000000000000000000000000011110",     --20
									 "0111100000000000000000000000000000011110",--1
								    "0111100000000000000000000000000000011110",--2
								    "0111100000000000000000000000000000011110",--3
								    "0111100000000000000000000000000000011110",--4
									 "0111100000000000000000000000000000011110",--5
									 "0111100000000000000000000000000000011110",--6
									 "0111100000000000000000000000000000011110",--7
									 "0111100000000000000000000000000000011110",--8
									 "0111100000000000000000000000000000011110",--9
								    "0111100000000000000000000000000000011110",--10         
								    "0111100000000000000000000000000000011110",--11
								    "0111100000000000000000000000000000011110",--12
								    "0111100000000000000000000000000000011110",--13
								    "0111100000000000000000000000000000011110",--14
								    "0111100000000000000000000000000000011110",--15
								    "0111100000000000000000000000000000011110",--16
								    "0111100000000000000000000000000000011110",--17
								    "0111100000000000000000000000000000011110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0111111111111111111111111111111111111110",     --40
									 "0111111111111111111111111111111111111110",--1
								    "0111111111111111111111111111111111111110",--2
								    "0000000000000000000000000000000000011110",--3
								    "0000000000000000000000000000000000011110",--4
									 "0000000000000000000000000000000000011110",--5
									 "0000000000000000000000000000000000011110",--6
									 "0000000000000000000000000000000000011110",--7
									 "0000000000000000000000000000000000011110",--8
									 "0000000000000000000000000000000000011110",--9
								    "0000000000000000000000000000000000011110",--10         
								    "0000000000000000000000000000000000011110",--11
								    "0000000000000000000000000000000000011110",--12
								    "0000000000000000000000000000000000011110",--13
								    "0000000000000000000000000000000000011110",--14
								    "0000000000000000000000000000000000011110",--15
								    "0000000000000000000000000000000000011110",--16
								    "0000000000000000000000000000000000011110",--17
								    "0000000000000000000000000000000000011110",--18
								    "0000000000000000000000000000000000011110",--19
								    "0000000000000000000000000000000000011110",    --60
									 "0000000000000000000000000000000000011110",--1
								    "0000000000000000000000000000000000011110",--2
								    "0000000000000000000000000000000000011110",--3
								    "0000000000000000000000000000000000011110",--4
									 "0000000000000000000000000000000000011110",--5
									 "0000000000000000000000000000000000011110",--6
									 "0000000000000000000000000000000000011110",--7
									 "0000000000000000000000000000000000011110",--8
									 "0000000000000000000000000000000000011110",--9
								    "0000000000000000000000000000000000011110",--10         
								    "0000000000000000000000000000000000011110",--11
								    "0000000000000000000000000000000000011110",--12
								    "0000000000000000000000000000000000011110",--13
								    "0000000000000000000000000000000000011110",--14
								    "0000000000000000000000000000000000011110",--15
								    "0000000000000000000000000000000000011110",--16
								    "0000000000000000000000000000000000011110",--17
								    "0000000000000000000000000000000000011110",--18
								    "0000000000000000000000000000000000011110",--19
								    "0000000000000000000000000000000000000000");  --80
									 
									 
									 
      constant BM_5: HFZ :=("0000000000000000000000000000000000000000",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0111111111111111111111111111111111111110",--5
									 "0111100000000000000000000000000000000000",--6
									 "0111100000000000000000000000000000000000",--7
									 "0111100000000000000000000000000000000000",--8
									 "0111100000000000000000000000000000000000",--9
								    "0111100000000000000000000000000000000000",--10         --22222222222
								    "0111100000000000000000000000000000000000",--11                  --222222222222
								    "0111100000000000000000000000000000000000",--12
								    "0111100000000000000000000000000000000000",--13
								    "0111100000000000000000000000000000000000",--14
								    "0111100000000000000000000000000000000000",--15
								    "0111100000000000000000000000000000000000",--16
								    "0111100000000000000000000000000000000000",--17
								    "0111100000000000000000000000000000000000",--18
								    "0111100000000000000000000000000000000000",--19
								    "0111100000000000000000000000000000000000",     --20
									 "0111100000000000000000000000000000000000",--1
								    "0111100000000000000000000000000000000000",--2
								    "0111100000000000000000000000000000000000",--3
								    "0111100000000000000000000000000000000000",--4
									 "0111100000000000000000000000000000000000",--5
									 "0111100000000000000000000000000000000000",--6
									 "0111100000000000000000000000000000000000",--7
									 "0111100000000000000000000000000000000000",--8
									 "0111100000000000000000000000000000000000",--9
								    "0111100000000000000000000000000000000000",--10         
								    "0111100000000000000000000000000000000000",--11
								    "0111100000000000000000000000000000000000",--12
								    "0111100000000000000000000000000000000000",--13
								    "0111100000000000000000000000000000000000",--14
								    "0111100000000000000000000000000000000000",--15
								    "0111100000000000000000000000000000000000",--16
								    "0111100000000000000000000000000000000000",--17
								    "0111100000000000000000000000000000000000",--18
								    "0111111111111111111111111111111111111110",--19
								    "0111111111111111111111111111111111111110",     --40
									 "0111111111111111111111111111111111111110",--1
								    "0111111111111111111111111111111111111110",--2
								    "0000000000000000000000000000000000011110",--3
								    "0000000000000000000000000000000000011110",--4
									 "0000000000000000000000000000000000011110",--5
									 "0000000000000000000000000000000000011110",--6
									 "0000000000000000000000000000000000011110",--7
									 "0000000000000000000000000000000000011110",--8
									 "0000000000000000000000000000000000011110",--9
								    "0000000000000000000000000000000000011110",--10         
								    "0000000000000000000000000000000000011110",--11
								    "0000000000000000000000000000000000011110",--12
								    "0000000000000000000000000000000000011110",--13
								    "0000000000000000000000000000000000011110",--14
								    "0000000000000000000000000000000000011110",--15
								    "0000000000000000000000000000000000011110",--16
								    "0000000000000000000000000000000000011110",--17
								    "0000000000000000000000000000000000011110",--18
								    "0000000000000000000000000000000000011110",--19
								    "0000000000000000000000000000000000011110",    --60
									 "0000000000000000000000000000000000011110",--1
								    "0000000000000000000000000000000000011110",--2
								    "0000000000000000000000000000000000011110",--3
								    "0000000000000000000000000000000000011110",--4
									 "0000000000000000000000000000000000011110",--5
									 "0000000000000000000000000000000000011110",--6
									 "0000000000000000000000000000000000011110",--7
									 "0000000000000000000000000000000000011110",--8
									 "0000000000000000000000000000000000011110",--9
								    "0000000000000000000000000000000000011110",--10         
								    "0000000000000000000000000000000000011110",--11
								    "0000000000000000000000000000000000011110",--12
								    "0000000000000000000000000000000000011110",--13
								    "0000000000000000000000000000000000011110",--14
								    "0000000000000000000000000000000000011110",--15
								    "0111111111111111111111111111111111111110",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0000000000000000000000000000000000000000");  --80
									 
									 
      constant BM_6: HFZ :=("0000000000000000000000000000000000000000",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0111111111111111111111111111111111111110",--5
									 "0111100000000000000000000000000000000000",--6
									 "0111100000000000000000000000000000000000",--7
									 "0111100000000000000000000000000000000000",--8
									 "0111100000000000000000000000000000000000",--9
								    "0111100000000000000000000000000000000000",--10         --22222222222
								    "0111100000000000000000000000000000000000",--11                  --222222222222
								    "0111100000000000000000000000000000000000",--12
								    "0111100000000000000000000000000000000000",--13
								    "0111100000000000000000000000000000000000",--14
								    "0111100000000000000000000000000000000000",--15
								    "0111100000000000000000000000000000000000",--16
								    "0111100000000000000000000000000000000000",--17
								    "0111100000000000000000000000000000000000",--18
								    "0111100000000000000000000000000000000000",--19
								    "0111100000000000000000000000000000000000",     --20
									 "0111100000000000000000000000000000000000",--1
								    "0111100000000000000000000000000000000000",--2
								    "0111100000000000000000000000000000000000",--3
								    "0111100000000000000000000000000000000000",--4
									 "0111100000000000000000000000000000000000",--5
									 "0111100000000000000000000000000000000000",--6
									 "0111100000000000000000000000000000000000",--7
									 "0111100000000000000000000000000000000000",--8
									 "0111100000000000000000000000000000000000",--9
								    "0111100000000000000000000000000000000000",--10         
								    "0111100000000000000000000000000000000000",--11
								    "0111100000000000000000000000000000000000",--12
								    "0111100000000000000000000000000000000000",--13
								    "0111100000000000000000000000000000000000",--14
								    "0111100000000000000000000000000000000000",--15
								    "0111100000000000000000000000000000000000",--16
								    "0111100000000000000000000000000000000000",--17
								    "0111100000000000000000000000000000000000",--18
								    "0111111111111111111111111111111111111110",--19
								    "0111111111111111111111111111111111111110",     --40
									 "0111111111111111111111111111111111111110",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111100000000000000000000000000000011110",--3
								    "0111100000000000000000000000000000011110",--4
									 "0111100000000000000000000000000000011110",--5
									 "0111100000000000000000000000000000011110",--6
									 "0111100000000000000000000000000000011110",--7
									 "0111100000000000000000000000000000011110",--8
									 "0111100000000000000000000000000000011110",--9
								    "0111100000000000000000000000000000011110",--10         
								    "0111100000000000000000000000000000011110",--11
								    "0111100000000000000000000000000000011110",--12
								    "0111100000000000000000000000000000011110",--13
								    "0111100000000000000000000000000000011110",--14
								    "0111100000000000000000000000000000011110",--15
								    "0111100000000000000000000000000000011110",--16
								    "0111100000000000000000000000000000011110",--17
								    "0111100000000000000000000000000000011110",--18
								    "0111100000000000000000000000000000011110",--19
								    "0111100000000000000000000000000000011110",    --60
									 "0111100000000000000000000000000000011110",--1
								    "0111100000000000000000000000000000011110",--2
								    "0111100000000000000000000000000000011110",--3
								    "0111100000000000000000000000000000011110",--4
									 "0111100000000000000000000000000000011110",--5
									 "0111100000000000000000000000000000011110",--6
									 "0111100000000000000000000000000000011110",--7
									 "0111100000000000000000000000000000011110",--8
									 "0111100000000000000000000000000000011110",--9
								    "0111100000000000000000000000000000011110",--10         
								    "0111100000000000000000000000000000011110",--11
								    "0111100000000000000000000000000000011110",--12
								    "0111100000000000000000000000000000011110",--13
								    "0111100000000000000000000000000000011110",--14
								    "0111100000000000000000000000000000011110",--15
								    "0111111111111111111111111111111111111110",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0000000000000000000000000000000000000000");  --80
									 
									 
	   constant BM_7: HFZ :=("0000000000000000000000000000000000000000",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0111111111111111111111111111111111111110",--5
									 "0000000000000000000000000000000000011110",--6
									 "0000000000000000000000000000000000011110",--7
									 "0000000000000000000000000000000000011110",--8
									 "0000000000000000000000000000000000011110",--9
								    "0000000000000000000000000000000000011110",--10         --33333333
								    "0000000000000000000000000000000000011110",--11                
								    "0000000000000000000000000000000000011110",--12
								    "0000000000000000000000000000000000011110",--13
								    "0000000000000000000000000000000000011110",--14
								    "0000000000000000000000000000000000011110",--15
								    "0000000000000000000000000000000000011110",--16
								    "0000000000000000000000000000000000011110",--17
								    "0000000000000000000000000000000000011110",--18
								    "0000000000000000000000000000000000011110",--19
								    "0000000000000000000000000000000000011110",     --20
									 "0000000000000000000000000000000000011110",--1
								    "0000000000000000000000000000000000011110",--2
								    "0000000000000000000000000000000000011110",--3
								    "0000000000000000000000000000000000011110",--4
									 "0000000000000000000000000000000000011110",--5
									 "0000000000000000000000000000000000011110",--6
									 "0000000000000000000000000000000000011110",--7
									 "0000000000000000000000000000000000011110",--8
									 "0000000000000000000000000000000000011110",--9
								    "0000000000000000000000000000000000011110",--10         
								    "0000000000000000000000000000000000011110",--11
								    "0000000000000000000000000000000000011110",--12
								    "0000000000000000000000000000000000011110",--13
								    "0000000000000000000000000000000000011110",--14
								    "0000000000000000000000000000000000011110",--15
								    "0000000000000000000000000000000000011110",--16
								    "0000000000000000000000000000000000011110",--17
								    "0000000000000000000000000000000000011110",--18
								    "0000000000000000000000000000000000011110",--19
								    "0000000000000000000000000000000000011110",     --40
									 "0000000000000000000000000000000000011110",--1
								    "0000000000000000000000000000000000011110",--2
								    "0000000000000000000000000000000000011110",--3
								    "0000000000000000000000000000000000011110",--4
									 "0000000000000000000000000000000000011110",--5
									 "0000000000000000000000000000000000011110",--6
									 "0000000000000000000000000000000000011110",--7
									 "0000000000000000000000000000000000011110",--8
									 "0000000000000000000000000000000000011110",--9
								    "0000000000000000000000000000000000011110",--10         
								    "0000000000000000000000000000000000011110",--11
								    "0000000000000000000000000000000000011110",--12
								    "0000000000000000000000000000000000011110",--13
								    "0000000000000000000000000000000000011110",--14
								    "0000000000000000000000000000000000011110",--15
								    "0000000000000000000000000000000000011110",--16
								    "0000000000000000000000000000000000011110",--17
								    "0000000000000000000000000000000000011110",--18
								    "0000000000000000000000000000000000011110",--19
								    "0000000000000000000000000000000000011110",    --60
									 "0000000000000000000000000000000000011110",--1
								    "0000000000000000000000000000000000011110",--2
								    "0000000000000000000000000000000000011110",--3
								    "0000000000000000000000000000000000011110",--4
									 "0000000000000000000000000000000000011110",--5
									 "0000000000000000000000000000000000011110",--6
									 "0000000000000000000000000000000000011110",--7
									 "0000000000000000000000000000000000011110",--8
									 "0000000000000000000000000000000000011110",--9
								    "0000000000000000000000000000000000011110",--10         
								    "0000000000000000000000000000000000011110",--11
								    "0000000000000000000000000000000000011110",--12
								    "0000000000000000000000000000000000011110",--13
								    "0000000000000000000000000000000000011110",--14
								    "0000000000000000000000000000000000011110",--15
								    "0000000000000000000000000000000000011110",--16
								    "0000000000000000000000000000000000011110",--17
								    "0000000000000000000000000000000000011110",--18
								    "0000000000000000000000000000000000011110",--19
								    "0000000000000000000000000000000000000000");  --80
									 
	   constant BM_8: HFZ :=("0000000000000000000000000000000000000000",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0111111111111111111111111111111111111110",--5
									 "0111100000000000000000000000000000011110",--6
									 "0111100000000000000000000000000000011110",--7
									 "0111100000000000000000000000000000011110",--8
									 "0111100000000000000000000000000000011110",--9
								    "0111100000000000000000000000000000011110",--10         --22222222222
								    "0111100000000000000000000000000000011110",--11                  --222222222222
								    "0111100000000000000000000000000000011110",--12
								    "0111100000000000000000000000000000011110",--13
								    "0111100000000000000000000000000000011110",--14
								    "0111100000000000000000000000000000011110",--15
								    "0111100000000000000000000000000000011110",--16
								    "0111100000000000000000000000000000011110",--17
								    "0111100000000000000000000000000000011110",--18
								    "0111100000000000000000000000000000011110",--19
								    "0111100000000000000000000000000000011110",     --20
									 "0111100000000000000000000000000000011110",--1
								    "0111100000000000000000000000000000011110",--2
								    "0111100000000000000000000000000000011110",--3
								    "0111100000000000000000000000000000011110",--4
									 "0111100000000000000000000000000000011110",--5
									 "0111100000000000000000000000000000011110",--6
									 "0111100000000000000000000000000000011110",--7
									 "0111100000000000000000000000000000011110",--8
									 "0111100000000000000000000000000000011110",--9
								    "0111100000000000000000000000000000011110",--10         
								    "0111100000000000000000000000000000011110",--11
								    "0111100000000000000000000000000000011110",--12
								    "0111100000000000000000000000000000011110",--13
								    "0111100000000000000000000000000000011110",--14
								    "0111100000000000000000000000000000011110",--15
								    "0111100000000000000000000000000000011110",--16
								    "0111100000000000000000000000000000011110",--17
								    "0111100000000000000000000000000000011110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0111111111111111111111111111111111111110",     --40
									 "0111111111111111111111111111111111111110",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111100000000000000000000000000000011110",--3
								    "0111100000000000000000000000000000011110",--4
									 "0111100000000000000000000000000000011110",--5
									 "0111100000000000000000000000000000011110",--6
									 "0111100000000000000000000000000000011110",--7
									 "0111100000000000000000000000000000011110",--8
									 "0111100000000000000000000000000000011110",--9
								    "0111100000000000000000000000000000011110",--10         
								    "0111100000000000000000000000000000011110",--11
								    "0111100000000000000000000000000000011110",--12
								    "0111100000000000000000000000000000011110",--13
								    "0111100000000000000000000000000000011110",--14
								    "0111100000000000000000000000000000011110",--15
								    "0111100000000000000000000000000000011110",--16
								    "0111100000000000000000000000000000011110",--17
								    "0111100000000000000000000000000000011110",--18
								    "0111100000000000000000000000000000011110",--19
								    "0111100000000000000000000000000000011110",    --60
									 "0111100000000000000000000000000000011110",--1
								    "0111100000000000000000000000000000011110",--2
								    "0111100000000000000000000000000000011110",--3
								    "0111100000000000000000000000000000011110",--4
									 "0111100000000000000000000000000000011110",--5
									 "0111100000000000000000000000000000011110",--6
									 "0111100000000000000000000000000000011110",--7
									 "0111100000000000000000000000000000011110",--8
									 "0111100000000000000000000000000000011110",--9
								    "0111100000000000000000000000000000011110",--10         
								    "0111100000000000000000000000000000011110",--11
								    "0111100000000000000000000000000000011110",--12
								    "0111100000000000000000000000000000011110",--13
								    "0111100000000000000000000000000000011110",--14
								    "0111100000000000000000000000000000011110",--15
								    "0111111111111111111111111111111111111110",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0000000000000000000000000000000000000000");  --80
									 
									 
	   constant BM_9: HFZ :=("0000000000000000000000000000000000000000",--1
								    "0111111111111111111111111111111111111110",--2
								    "0111111111111111111111111111111111111110",--3
								    "0111111111111111111111111111111111111110",--4
									 "0111111111111111111111111111111111111110",--5
									 "0111100000000000000000000000000000011110",--6
									 "0111100000000000000000000000000000011110",--7
									 "0111100000000000000000000000000000011110",--8
									 "0111100000000000000000000000000000011110",--9
								    "0111100000000000000000000000000000011110",--10         --22222222222
								    "0111100000000000000000000000000000011110",--11                  --222222222222
								    "0111100000000000000000000000000000011110",--12
								    "0111100000000000000000000000000000011110",--13
								    "0111100000000000000000000000000000011110",--14
								    "0111100000000000000000000000000000011110",--15
								    "0111100000000000000000000000000000011110",--16
								    "0111100000000000000000000000000000011110",--17
								    "0111100000000000000000000000000000011110",--18
								    "0111100000000000000000000000000000011110",--19
								    "0111100000000000000000000000000000011110",     --20
									 "0111100000000000000000000000000000011110",--1
								    "0111100000000000000000000000000000011110",--2
								    "0111100000000000000000000000000000011110",--3
								    "0111100000000000000000000000000000011110",--4
									 "0111100000000000000000000000000000011110",--5
									 "0111100000000000000000000000000000011110",--6
									 "0111100000000000000000000000000000011110",--7
									 "0111100000000000000000000000000000011110",--8
									 "0111100000000000000000000000000000011110",--9
								    "0111100000000000000000000000000000011110",--10         
								    "0111100000000000000000000000000000011110",--11
								    "0111100000000000000000000000000000011110",--12
								    "0111100000000000000000000000000000011110",--13
								    "0111100000000000000000000000000000011110",--14
								    "0111100000000000000000000000000000011110",--15
								    "0111100000000000000000000000000000011110",--16
								    "0111100000000000000000000000000000011110",--17
								    "0111100000000000000000000000000000011110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0111111111111111111111111111111111111110",     --40
									 "0111111111111111111111111111111111111110",--1
								    "0111111111111111111111111111111111111110",--2
								    "0000000000000000000000000000000000011110",--3
								    "0000000000000000000000000000000000011110",--4
									 "0000000000000000000000000000000000011110",--5
									 "0000000000000000000000000000000000011110",--6
									 "0000000000000000000000000000000000011110",--7
									 "0000000000000000000000000000000000011110",--8
									 "0000000000000000000000000000000000011110",--9
								    "0000000000000000000000000000000000011110",--10         
								    "0000000000000000000000000000000000011110",--11
								    "0000000000000000000000000000000000011110",--12
								    "0000000000000000000000000000000000011110",--13
								    "0000000000000000000000000000000000011110",--14
								    "0000000000000000000000000000000000011110",--15
								    "0000000000000000000000000000000000011110",--16
								    "0000000000000000000000000000000000011110",--17
								    "0000000000000000000000000000000000011110",--18
								    "0000000000000000000000000000000000011110",--19
								    "0000000000000000000000000000000000011110",    --60
									 "0000000000000000000000000000000000011110",--1
								    "0000000000000000000000000000000000011110",--2
								    "0000000000000000000000000000000000011110",--3
								    "0000000000000000000000000000000000011110",--4
									 "0000000000000000000000000000000000011110",--5
									 "0000000000000000000000000000000000011110",--6
									 "0000000000000000000000000000000000011110",--7
									 "0000000000000000000000000000000000011110",--8
									 "0000000000000000000000000000000000011110",--9
								    "0000000000000000000000000000000000011110",--10         
								    "0000000000000000000000000000000000011110",--11
								    "0000000000000000000000000000000000011110",--12
								    "0000000000000000000000000000000000011110",--13
								    "0000000000000000000000000000000000011110",--14
								    "0000000000000000000000000000000000011110",--15
								    "0111111111111111111111111111111111111110",--16
								    "0111111111111111111111111111111111111110",--17
								    "0111111111111111111111111111111111111110",--18
								    "0111111111111111111111111111111111111110",--19
								    "0000000000000000000000000000000000000000");  --80
									 

								

									 
	
constant BM_iki_nokta:HFZ:=("0000000000000000000000000000000000000000",--1
								    "0000000000000000000000000000000000000000",--2
								    "0000000000000000000000000000000000000000",--3
								    "0000000000000000000000000000000000000000",--4
									 "0000000000000000000000000000000000000000",--5
									 "0000000000000000000000000000000000000000",--6
									 "0000000000000000000000000000000000000000",--7
									 "0000000000000000000000000000000000000000",--8
									 "0000000000000000000000000000000000000000",--9
								    "0000000000000000000000000000000000000000",--10         --BOS
								    "0000000000000000000000000000000000000000",--11
								    "0000000000000000000000000000000000000000",--12
								    "0000000000000000000000000000000000000000",--13
								    "0000000000000000000000000000000000000000",--14
								    "0000000000111111111111111111110000000000",--15
								    "0000000000111111111111111111110000000000",--16
								    "0000000000111111111111111111110000000000",--17
								    "0000000000111111111111111111110000000000",--18
								    "0000000000111111111111111111110000000000",--19
								    "0000000000111111111111111111110000000000",     --20
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000111111111111111111110000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000",
									 "0000000000000000000000000000000000000000");

begin
	--get 40Mhz clock
	c1_pll2: PLL port map(clk_in_clk=>CLOCK_50 , reset_reset=>reset , clk_out_clk=>clk_40);
	
	clk_divider: process(CLOCK_50)
	begin
		if rising_edge(CLOCK_50) then
			clk_div <= clk_div + 1;
		end if;
	end process;
	clk15 <= clk_div(15);
	
	
	--get 1Hz clock
	process(CLOCK_50)
	variable cnt : integer;
   begin
		if rising_edge(CLOCK_50) then
			if SW(1) = '0' then
				 if (cnt<10000000) then
					 cnt:=cnt+1;
				 else
					 clk_1hz <= NOT(clk_1hz);
					 cnt:=0;
			    end if;
			else
				if (cnt=24999999) then
					 clk_1hz <= NOT(clk_1hz);
					 cnt:=0;
				 else
               cnt:=cnt+1;
			    end if;
			end if;
     end if;
	end process;
	

	--0 to 59 counter
	process(clk_1hz,SW(0),KEY(0),KEY(1),clk15) 
	begin
		if rst = '0' then
			cntr59 <= 0;
			cntr59_min <= 0;
			cntr59_hour <= 0;
		elsif rising_edge(clk_1hz) then
			if SW(0) = '1' then
				if enable = '1' then
					if cntr59 > 0 then
						cntr59 <= cntr59  - 1;
					else
						cntr59 <= 59;
						cntr59_min <= cntr59_min - 1;
						if cntr59_min = 0 then
							cntr59_min <= 59;
							cntr59_hour <= cntr59_hour - 1;
							if cntr59_hour = 0 then
								cntr59_hour <= 0;
								cntr59_min <= 0;
								cntr59 <= 0;
								enable <= '0';
								GPIO_0(0) <= '1';
							end if;
						end if;
					end if;
				end if;
			else
				if KEY(0)='0' then
					enable <= '1';
					GPIO_0(0) <= '0';
					if cntr59 < 59 then
						cntr59 <= cntr59  + 1;
					else
						cntr59 <= 0;
					end if;
						
				elsif KEY(1)='0' then
					enable <= '1';
					GPIO_0(0) <= '0';
					cntr59_min <= cntr59_min+1;
					if cntr59_min = 59 then
						cntr59_min <= 0;
					end if;
					
				elsif KEY(2)='0' then
					cntr59_hour <= cntr59_hour+1;
					if cntr59_hour = 59 then
						cntr59_hour <= 0;
					end if;
				end if;
			end if;
		end if;	
	end process;
	
-------------------------------------------
	VGA_CLK<=clk_40;
	VGA_BLANK <= (VGA_HS and VGA_VS);
-------------------------------------------
	
Horizontal_position_counter:process(clk_40)
begin
	if(clk_40'event and clk_40 = '1')then
		if (hPos = (HD + HFP + HSP + HBP)) then
			hPos <= 0;
		else
			hPos <= hPos + 1;
		end if;
	end if;
end process;


Vertical_position_counter:process(clk_40, hPos)
begin
	if(clk_40'event and clk_40 = '1')then
		if(hPos = (HD + HFP + HSP + HBP))then
			if (vPos = (VD + VFP + VSP + VBP)) then
				vPos <= 0;
			else
				vPos <= vPos + 1;
			end if;
		end if;
	end if;
end process;
	
Horizontal_Synchronisation:process(clk_40, hPos)
begin
	if(clk_40'event and clk_40 = '1')then
		if((hPos <= (HD + HFP)) OR (hPos > HD + HFP + HSP))then
			VGA_HS <= '1';
		else
			VGA_HS <= '0';
		end if;
	end if;
end process;


Vertical_Synchronisation:process(clk_40, vPos)
begin
	if(clk_40'event and clk_40 = '1')then
		if((vPos <= (VD + VFP)) OR (vPos > VD + VFP + VSP))then
			VGA_VS <= '1';
		else
			VGA_VS <= '0';
		end if;
	end if;
end process;


video_on:process(clk_40, hPos, vPos)
begin
	if(clk_40'event and clk_40 = '1')then
		if(hPos <= HD and vPos <= VD)then
			videoOn <= '1';
		else
			videoOn <= '0';
		end if;
	end if;
end process;
	
draw:process(clk_40, clk_1hz, hPos, vPos, videoOn)
variable bmbit: std_logic;
variable bmbit1: std_logic;
variable bmbit2: std_logic;
variable bmbit3: std_logic;
variable bmbit4: std_logic;
variable bmbit5: std_logic;
variable bmbit6: std_logic;
variable bmbit7: std_logic;
variable bmbit8: std_logic;
begin
	if(clk_40'event and clk_40 = '1')then
		if(videoOn = '1')then
			if ((hpos>=100 AND hpos<200) AND (vpos>100 AND vpos<200)) THEN
				VGA_R <= "1111111111";
				VGA_G <= "1111111111";
				VGA_B <= "0000000000";
			else
				VGA_R <= "0000000000";
				VGA_G <= "0000000000";
				VGA_B <= "0000000000";
			end if;
			
		
			
			if(cntr59 mod 10 = 0) then	
				bmbit:= BM_0(vpos mod 80)(hpos mod 40);
			elsif(cntr59 mod 10 = 1) then	
				bmbit:= BM_1(vpos mod 80)(hpos mod 40);	
			elsif(cntr59 mod 10 = 2) then	
				bmbit:= BM_2(vpos mod 80)(hpos mod 40);
			elsif(cntr59 mod 10 = 3) then	
				bmbit:= BM_3(vpos mod 80)(hpos mod 40);
			elsif(cntr59 mod 10 = 4) then	
				bmbit:= BM_4(vpos mod 80)(hpos mod 40);
			elsif(cntr59 mod 10 = 5) then	
				bmbit:= BM_5(vpos mod 80)(hpos mod 40);
			elsif(cntr59 mod 10 = 6) then	
				bmbit:= BM_6(vpos mod 80)(hpos mod 40);
			elsif(cntr59 mod 10 = 7) then	
				bmbit:= BM_7(vpos mod 80)(hpos mod 40);
			elsif(cntr59 mod 10 = 8) then	
				bmbit:= BM_8(vpos mod 80)(hpos mod 40);
			elsif(cntr59 mod 10 = 9) then	
				bmbit:= BM_9(vpos mod 80)(hpos mod 40);
			end if;
			

			if cntr59 < 10 then 
				bmbit2:= BM_0(vpos mod 80)(hpos mod 40);
			elsif cntr59 < 20 then 
				bmbit2:=BM_1(vpos mod 80)(hpos mod 40);
			elsif cntr59 < 30 then  
				bmbit2:= BM_2(vpos mod 80)(hpos mod 40);
			elsif cntr59 < 40 then 
				bmbit2:= BM_3(vpos mod 80)(hpos mod 40);
			elsif cntr59 < 50 then  
				bmbit2:= BM_4(vpos mod 80)(hpos mod 40);
			elsif cntr59 <60 then  
				bmbit2:= BM_5(vpos mod 80)(hpos mod 40);
			elsif cntr59 =60 then  
				bmbit2:= BM_0(vpos mod 80)(hpos mod 40);
			end if;
			
			
			--dakika için
			if(cntr59_min mod 10 = 0) then	
				bmbit4:= BM_0(vpos mod 80)(hpos mod 40);
			elsif(cntr59_min mod 10 = 1) then	
				bmbit4:= BM_1(vpos mod 80)(hpos mod 40);	
			elsif(cntr59_min mod 10 = 2) then	
				bmbit4:= BM_2(vpos mod 80)(hpos mod 40);
			elsif(cntr59_min mod 10 = 3) then	
				bmbit4:= BM_3(vpos mod 80)(hpos mod 40);
			elsif(cntr59_min mod 10 = 4) then	
				bmbit4:= BM_4(vpos mod 80)(hpos mod 40);
			elsif(cntr59_min mod 10 = 5) then	
				bmbit4:= BM_5(vpos mod 80)(hpos mod 40);
			elsif(cntr59_min mod 10 = 6) then	
				bmbit4:= BM_6(vpos mod 80)(hpos mod 40);
			elsif(cntr59_min mod 10 = 7) then	
				bmbit4:= BM_7(vpos mod 80)(hpos mod 40);
			elsif(cntr59_min mod 10 = 8) then	
				bmbit4:= BM_8(vpos mod 80)(hpos mod 40);
			elsif(cntr59_min mod 10 = 9) then	
				bmbit4:= BM_9(vpos mod 80)(hpos mod 40);
			end if;
			
			if cntr59_min < 10 then 
				bmbit5:= BM_0(vpos mod 80)(hpos mod 40);
			elsif cntr59_min < 20 then 
				bmbit5:=BM_1(vpos mod 80)(hpos mod 40);
			elsif cntr59_min < 30 then  
				bmbit5:= BM_2(vpos mod 80)(hpos mod 40);
			elsif cntr59_min < 40 then 
				bmbit5:= BM_3(vpos mod 80)(hpos mod 40);
			elsif cntr59_min < 50 then  
				bmbit5:= BM_4(vpos mod 80)(hpos mod 40);
			elsif cntr59_min <60 then  
				bmbit5:= BM_5(vpos mod 80)(hpos mod 40);
			elsif cntr59_min =60 then  
				bmbit5:= BM_0(vpos mod 80)(hpos mod 40);
			end if;
			
			
			
			--saat için
			if(cntr59_hour mod 10 = 0) then	
				bmbit6:= BM_0(vpos mod 80)(hpos mod 40);
			elsif(cntr59_hour mod 10 = 1) then	
				bmbit6:= BM_1(vpos mod 80)(hpos mod 40);	
			elsif(cntr59_hour mod 10 = 2) then	
				bmbit6:= BM_2(vpos mod 80)(hpos mod 40);
			elsif(cntr59_hour mod 10 = 3) then	
				bmbit6:= BM_3(vpos mod 80)(hpos mod 40);
			elsif(cntr59_hour mod 10 = 4) then	
				bmbit6:= BM_4(vpos mod 80)(hpos mod 40);
			elsif(cntr59_hour mod 10 = 5) then	
				bmbit6:= BM_5(vpos mod 80)(hpos mod 40);
			elsif(cntr59_hour mod 10 = 6) then	
				bmbit6:= BM_6(vpos mod 80)(hpos mod 40);
			elsif(cntr59_hour mod 10 = 7) then	
				bmbit6:= BM_7(vpos mod 80)(hpos mod 40);
			elsif(cntr59_hour mod 10 = 8) then	
				bmbit6:= BM_8(vpos mod 80)(hpos mod 40);
			elsif(cntr59_hour mod 10 = 9) then	
				bmbit6:= BM_9(vpos mod 80)(hpos mod 40);
			end if;
			
			if cntr59_hour < 10 then 
				bmbit7:= BM_0(vpos mod 80)(hpos mod 40);
			elsif cntr59_hour < 20 then 
				bmbit7:=BM_1(vpos mod 80)(hpos mod 40);
			elsif cntr59_hour < 30 then  
				bmbit7:= BM_2(vpos mod 80)(hpos mod 40);
			elsif cntr59_hour < 40 then 
				bmbit7:= BM_3(vpos mod 80)(hpos mod 40);
			elsif cntr59_hour < 50 then  
				bmbit7:= BM_4(vpos mod 80)(hpos mod 40);
			elsif cntr59_hour <60 then  
				bmbit7:= BM_5(vpos mod 80)(hpos mod 40);
			elsif cntr59_hour =60 then  
				bmbit7:= BM_0(vpos mod 80)(hpos mod 40);
			end if;
				
			if ((hpos>=200 AND hpos<240) AND (vpos>=320 AND vpos<400)) THEN
				if bmbit7='1' then
					VGA_R <= "1111111111";
					VGA_G <= "0000000000";
					VGA_B <= "0000000000";
				else	
					VGA_R <= "1111111111";
					VGA_G <= "1111111111";
					VGA_B <= "1111111111";
				end if;
			end if;
		
			if ((hpos>=240 AND hpos<280) AND (vpos>=320 AND vpos<400)) THEN
				if bmbit6='1' then
					VGA_R <= "1111111111";
					VGA_G <= "0000000000";
					VGA_B <= "0000000000";
				else	
					VGA_R <= "1111111111";
					VGA_G <= "1111111111";
					VGA_B <= "1111111111";
				end if;
			end if;
				
			if ((hpos>=280 AND hpos<320) AND (vpos>=320 AND vpos<400)) THEN
				bmbit8:= BM_iki_nokta(vpos mod 80)(hpos mod 40);
				if bmbit8='1' then
					VGA_R <= "1111111111";
					VGA_G <= "0000000000";
					VGA_B <= "0000000000";
				else	
					VGA_R <= "1111111111";
					VGA_G <= "1111111111";
					VGA_B <= "1111111111";
				end if;
			end if;
			
			if ((hpos>=320 AND hpos<360) AND (vpos>=320 AND vpos<400)) THEN
				if bmbit5='1' then
					VGA_R <= "1111111111";
					VGA_G <= "0000000000";
					VGA_B <= "0000000000";
				else	
					VGA_R <= "1111111111";
					VGA_G <= "1111111111";
					VGA_B <= "1111111111";
				end if;
			end if;
			
			if ((hpos>=360 AND hpos<400) AND (vpos>=320 AND vpos<400)) THEN
				if bmbit4='1' then
					VGA_R <= "1111111111";
					VGA_G <= "0000000000";
					VGA_B <= "0000000000";
				else	
					VGA_R <= "1111111111";
					VGA_G <= "1111111111";
					VGA_B <= "1111111111";
				end if;
			end if;
			
			--asagıdakiler saniye içindir.
			if ((hpos>=400 AND hpos<440) AND (vpos>=320 AND vpos<400)) THEN
				bmbit3:= BM_iki_nokta(vpos mod 80)(hpos mod 40);
				if bmbit3='1' then
					VGA_R <= "1111111111";
					VGA_G <= "0000000000";
					VGA_B <= "0000000000";
				else	
					VGA_R <= "1111111111";
					VGA_G <= "1111111111";
					VGA_B <= "1111111111";
				end if;
			end if;
			
			if ((hpos>=440 AND hpos<480) AND (vpos>=320 AND vpos<400)) THEN
				if bmbit2 = '1' then
					VGA_R <= "1111111111";
					VGA_G <= "0000000000";
					VGA_B <= "0000000000";
				else	
					VGA_R <= "1111111111";
					VGA_G <= "1111111111";
					VGA_B <= "1111111111";
				end if;
			end if;
			
		   if ((hpos>=480 AND hpos<520) AND (vpos>=320 AND vpos<400)) THEN
				if bmbit = '1' then
					VGA_R <= "1111111111";
					VGA_G <= "0000000000";
					VGA_B <= "0000000000";
				else	
					VGA_R <= "1111111111";
					VGA_G <= "1111111111";
					VGA_B <= "1111111111";
				end if;
			end if;
			

		else
			VGA_R <= "0000000000";
			VGA_G <= "0000000000";
			VGA_B <= "0000000000";
		end if;
	end if;
end process;

	
end architecture;
